module corebit_not (
    input in,
    output out
);
  assign out = ~in;
endmodule

