module Main (
    input [2:0] I0 [5:0][3:0],
    input I1__0,
    input [2:0] I1__1,
    output [2:0] O0 [1:0][3:0],
    output [2:0] O1 [3:0][3:0]
);
assign O0 = {{I0[1][1],I0[1][2],I0[1][3],I0[1][0]},{I0[0][1],I0[0][2],I0[0][3],I0[0][0]}};
assign O1 = {{{I0[5][1][1],I0[5][1][2],I0[5][1][0]},{I0[5][2][1],I0[5][2][2],I0[5][2][0]},{I0[5][3][1],I0[5][3][2],I0[5][3][0]},{I0[5][0][1],I0[5][0][2],I0[5][0][0]}},{{I0[4][1][1],I0[4][1][2],I0[4][1][0]},{I0[4][2][1],I0[4][2][2],I0[4][2][0]},{I0[4][3][1],I0[4][3][2],I0[4][3][0]},{I0[4][0][1],I0[4][0][2],I0[4][0][0]}},{{I0[3][1][1],I0[3][1][2],I0[3][1][0]},{I0[3][2][1],I0[3][2][2],I0[3][2][0]},{I0[3][3][1],I0[3][3][2],I0[3][3][0]},{I0[3][0][1],I0[3][0][2],I0[3][0][0]}},{{I0[2][1][1],I0[2][1][2],I0[2][1][0]},{I0[2][2][1],I0[2][2][2],I0[2][2][0]},{I0[2][3][1],I0[2][3][2],I0[2][3][0]},{I0[2][0][1],I0[2][0][2],I0[2][0][0]}}};
endmodule

