// Module `SB_RAM40_4K` defined externally
module top (
    input [15:0] MASK,
    input [10:0] RADDR,
    input RCLK,
    input RCLKE,
    output [15:0] RDATA,
    input RE,
    input [10:0] WADDR,
    input WCLK,
    input WCLKE,
    input [15:0] WDATA,
    input WE
);
wire [15:0] SB_RAM40_4K_inst0_RDATA;
wire [10:0] SB_RAM40_4K_inst0_RADDR;
wire SB_RAM40_4K_inst0_RCLK;
wire SB_RAM40_4K_inst0_RCLKE;
wire SB_RAM40_4K_inst0_RE;
wire SB_RAM40_4K_inst0_WCLK;
wire SB_RAM40_4K_inst0_WCLKE;
wire SB_RAM40_4K_inst0_WE;
wire [10:0] SB_RAM40_4K_inst0_WADDR;
wire [15:0] SB_RAM40_4K_inst0_MASK;
wire [15:0] SB_RAM40_4K_inst0_WDATA;
assign SB_RAM40_4K_inst0_RADDR = RADDR;
assign SB_RAM40_4K_inst0_RCLK = RCLK;
assign SB_RAM40_4K_inst0_RCLKE = RCLKE;
assign SB_RAM40_4K_inst0_RE = RE;
assign SB_RAM40_4K_inst0_WCLK = WCLK;
assign SB_RAM40_4K_inst0_WCLKE = WCLKE;
assign SB_RAM40_4K_inst0_WE = WE;
assign SB_RAM40_4K_inst0_WADDR = WADDR;
assign SB_RAM40_4K_inst0_MASK = MASK;
assign SB_RAM40_4K_inst0_WDATA = WDATA;
SB_RAM40_4K #(
    .INIT_0(256'h0000000000000000000000000000000000000000000000000000000000ff00fe),
    .INIT_1(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_8(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_9(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .READ_MODE(0),
    .WRITE_MODE(0)
) SB_RAM40_4K_inst0 (
    .RDATA(SB_RAM40_4K_inst0_RDATA),
    .RADDR(SB_RAM40_4K_inst0_RADDR),
    .RCLK(SB_RAM40_4K_inst0_RCLK),
    .RCLKE(SB_RAM40_4K_inst0_RCLKE),
    .RE(SB_RAM40_4K_inst0_RE),
    .WCLK(SB_RAM40_4K_inst0_WCLK),
    .WCLKE(SB_RAM40_4K_inst0_WCLKE),
    .WE(SB_RAM40_4K_inst0_WE),
    .WADDR(SB_RAM40_4K_inst0_WADDR),
    .MASK(SB_RAM40_4K_inst0_MASK),
    .WDATA(SB_RAM40_4K_inst0_WDATA)
);
assign RDATA = SB_RAM40_4K_inst0_RDATA;
endmodule

