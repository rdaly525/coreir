module Main (input [4:0] I, output [4:0] O);
wire [4:0] x;
assign x = I;
assign O = x;
endmodule

