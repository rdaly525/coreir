module Main (input I, output O);
wire x;
assign x = I;
assign O = x;
endmodule

